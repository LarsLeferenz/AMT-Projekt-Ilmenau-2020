-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Wed Mar 11 10:56:36 2020

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY fahrstrecke_einlesen IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        sl : OUT STD_LOGIC;
        sr : OUT STD_LOGIC;
        sk : OUT STD_LOGIC;
        dl : OUT STD_LOGIC;
        dr : OUT STD_LOGIC;
        st : OUT STD_LOGIC;
        y0 : OUT STD_LOGIC;
        y1 : OUT STD_LOGIC;
        y2 : OUT STD_LOGIC;
        y3 : OUT STD_LOGIC;
        triggerNext : OUT STD_LOGIC
    );
END fahrstrecke_einlesen;

ARCHITECTURE BEHAVIOR OF fahrstrecke_einlesen IS
    TYPE type_fstate IS (init);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset)
    BEGIN
        IF (reset='0') THEN
            reg_fstate <= init;
            sl <= '0';
            sr <= '0';
            sk <= '0';
            dl <= '0';
            dr <= '0';
            st <= '0';
            y0 <= '0';
            y1 <= '0';
            y2 <= '0';
            y3 <= '0';
            triggerNext <= '0';
        ELSE
            sl <= '0';
            sr <= '0';
            sk <= '0';
            dl <= '0';
            dr <= '0';
            st <= '0';
            y0 <= '0';
            y1 <= '0';
            y2 <= '0';
            y3 <= '0';
            triggerNext <= '0';
            CASE fstate IS
                WHEN init =>
                    reg_fstate <= init;

                    st <= '0';

                    triggerNext <= '0';

                    sk <= '0';

                    y3 <= '0';

                    sl <= '0';

                    sr <= '0';

                    dr <= '0';

                    y1 <= '0';

                    y2 <= '0';

                    y0 <= '0';

                    dl <= '0';
                WHEN OTHERS => 
                    sl <= 'X';
                    sr <= 'X';
                    sk <= 'X';
                    dl <= 'X';
                    dr <= 'X';
                    st <= 'X';
                    y0 <= 'X';
                    y1 <= 'X';
                    y2 <= 'X';
                    y3 <= 'X';
                    triggerNext <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
