-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Wed Aug 19 14:04:58 2020

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY vierbit_Save IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        write : IN STD_LOGIC := '0';
        x1 : IN STD_LOGIC := '0';
        x0 : IN STD_LOGIC := '0';
        read : IN STD_LOGIC := '0';
        y1 : OUT STD_LOGIC;
        y0 : OUT STD_LOGIC;
        y1arr : OUT STD_LOGIC;
        y0arr : OUT STD_LOGIC
    );
END vierbit_Save;

ARCHITECTURE BEHAVIOR OF vierbit_Save IS
    TYPE type_fstate IS (z0,z1,z2,z3);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,write,x1,x0,read)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= z0;
            y1 <= '0';
            y0 <= '0';
            y1arr <= '0';
            y0arr <= '0';
        ELSE
            y1 <= '0';
            y0 <= '0';
            y1arr <= '0';
            y0arr <= '0';
            CASE fstate IS
                WHEN z0 =>
                    IF ((((write = '1') AND (x0 = '1')) AND NOT((x1 = '1')))) THEN
                        reg_fstate <= z1;
                    ELSIF ((((write = '1') AND (x1 = '1')) AND NOT((x0 = '1')))) THEN
                        reg_fstate <= z2;
                    ELSIF ((((write = '1') AND (x0 = '1')) AND (x1 = '1'))) THEN
                        reg_fstate <= z3;
                    ELSIF ((NOT((write = '1')) OR (NOT((x0 = '1')) AND NOT((x1 = '1'))))) THEN
                        reg_fstate <= z0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= z0;
                    END IF;

                    y1 <= '0';

                    y0 <= '0';
                WHEN z1 =>
                    IF (((write = '1') AND (NOT((x0 = '1')) OR (x1 = '1')))) THEN
                        reg_fstate <= z0;
                    ELSIF ((NOT((write = '1')) OR ((x0 = '1') AND NOT((x1 = '1'))))) THEN
                        reg_fstate <= z1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= z1;
                    END IF;

                    y0arr <= '1';

                    y1 <= '0';

                    IF ((read = '1')) THEN
                        y0 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        y0 <= '0';
                    END IF;
                WHEN z2 =>
                    IF (((write = '1') AND (NOT((x1 = '1')) OR (x0 = '1')))) THEN
                        reg_fstate <= z0;
                    ELSIF ((NOT((write = '1')) OR (NOT((x0 = '1')) AND (x1 = '1')))) THEN
                        reg_fstate <= z2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= z2;
                    END IF;

                    y1arr <= '1';

                    IF ((read = '1')) THEN
                        y1 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        y1 <= '0';
                    END IF;

                    y0 <= '0';
                WHEN z3 =>
                    IF (((write = '1') AND (NOT((x0 = '1')) OR NOT((x1 = '1'))))) THEN
                        reg_fstate <= z0;
                    ELSIF ((NOT((write = '1')) OR ((x0 = '1') AND (x1 = '1')))) THEN
                        reg_fstate <= z3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= z3;
                    END IF;

                    y0arr <= '1';

                    y1arr <= '1';

                    IF ((read = '1')) THEN
                        y1 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        y1 <= '0';
                    END IF;

                    IF ((read = '1')) THEN
                        y0 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        y0 <= '0';
                    END IF;
                WHEN OTHERS => 
                    y1 <= 'X';
                    y0 <= 'X';
                    y1arr <= 'X';
                    y0arr <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
