-- Copyright (C) 2019  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 19.1.0 Build 670 09/22/2019 SJ Lite Edition
-- Created on Fri Aug 28 17:43:44 2020

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY HEX_zweiverschoben IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        x : IN STD_LOGIC := '0';
        x2 : IN STD_LOGIC := '0';
        b3 : OUT STD_LOGIC;
        b2 : OUT STD_LOGIC;
        b1 : OUT STD_LOGIC;
        b0 : OUT STD_LOGIC;
        y : OUT STD_LOGIC
    );
END HEX_zweiverschoben;

ARCHITECTURE BEHAVIOR OF HEX_zweiverschoben IS
    TYPE type_fstate IS (Z0,Z1,Z2,Z3,Z4,Z5,Z6,Z7,Z8,Z9,ZA,ZB,ZC,ZD,ZE,ZF,vor,vor2,vor3);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= vor;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,x,x2)
    BEGIN
        b3 <= '0';
        b2 <= '0';
        b1 <= '0';
        b0 <= '0';
        y <= '0';
        CASE fstate IS
            WHEN Z0 =>
                IF (NOT((x = '1'))) THEN
                    reg_fstate <= Z0;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= Z1;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z0;
                END IF;

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;
                y <= '1';

                b3 <= '0';

                b1 <= '0';

                b2 <= '0';

                b0 <= '0';
            WHEN Z1 =>
                IF (NOT((x2 = '1'))) THEN
                    reg_fstate <= Z1;
                ELSIF ((x2 = '1')) THEN
                    reg_fstate <= Z2;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z1;
                END IF;

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;

                b3 <= '0';

                b1 <= '0';

                b2 <= '0';

                b0 <= '1';
            WHEN Z2 =>
                IF (NOT((x = '1'))) THEN
                    reg_fstate <= Z2;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= Z3;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z2;
                END IF;

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;

                b3 <= '0';

                b1 <= '1';

                b2 <= '0';

                b0 <= '0';
            WHEN Z3 =>
                IF (NOT((x2 = '1'))) THEN
                    reg_fstate <= Z3;
                ELSIF ((x2 = '1')) THEN
                    reg_fstate <= Z4;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z3;
                END IF;

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;

                b3 <= '0';

                b1 <= '1';

                b2 <= '0';

                b0 <= '1';
            WHEN Z4 =>
                IF (NOT((x = '1'))) THEN
                    reg_fstate <= Z4;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= Z5;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z4;
                END IF;

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;

                b3 <= '0';

                b1 <= '0';

                b2 <= '1';

                b0 <= '0';
            WHEN Z5 =>
                IF (NOT((x2 = '1'))) THEN
                    reg_fstate <= Z5;
                ELSIF ((x2 = '1')) THEN
                    reg_fstate <= Z6;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z5;
                END IF;

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;

                b3 <= '0';

                b1 <= '0';

                b2 <= '1';

                b0 <= '1';
            WHEN Z6 =>
                IF (NOT((x = '1'))) THEN
                    reg_fstate <= Z6;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= Z7;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z6;
                END IF;

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;

                b3 <= '0';

                b1 <= '1';

                b2 <= '1';

                b0 <= '0';
            WHEN Z7 =>
                IF (NOT((x2 = '1'))) THEN
                    reg_fstate <= Z7;
                ELSIF ((x2 = '1')) THEN
                    reg_fstate <= Z8;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z7;
                END IF;

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;

                b3 <= '0';

                b1 <= '1';

                b2 <= '1';

                b0 <= '1';
            WHEN Z8 =>
                IF (NOT((x = '1'))) THEN
                    reg_fstate <= Z8;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= Z9;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z8;
                END IF;

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;

                b3 <= '1';

                b1 <= '0';

                b2 <= '0';

                b0 <= '0';
            WHEN Z9 =>
                IF (NOT((x2 = '1'))) THEN
                    reg_fstate <= Z9;
                ELSIF ((x2 = '1')) THEN
                    reg_fstate <= ZA;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z9;
                END IF;

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;

                b3 <= '1';

                b1 <= '0';

                b2 <= '0';

                b0 <= '1';
            WHEN ZA =>
                IF (NOT((x = '1'))) THEN
                    reg_fstate <= ZA;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= ZB;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= ZA;
                END IF;

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;

                b3 <= '1';

                b1 <= '1';

                b2 <= '0';

                b0 <= '0';
            WHEN ZB =>
                IF (NOT((x2 = '1'))) THEN
                    reg_fstate <= ZB;
                ELSIF ((x2 = '1')) THEN
                    reg_fstate <= ZC;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= ZB;
                END IF;

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;

                b3 <= '1';

                b1 <= '1';

                b2 <= '0';

                b0 <= '1';
            WHEN ZC =>
                IF (NOT((x = '1'))) THEN
                    reg_fstate <= ZC;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= ZD;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= ZC;
                END IF;

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;

                b3 <= '1';

                b1 <= '0';

                b2 <= '1';

                b0 <= '0';
            WHEN ZD =>
                IF (NOT((x2 = '1'))) THEN
                    reg_fstate <= ZD;
                ELSIF ((x2 = '1')) THEN
                    reg_fstate <= ZE;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= ZD;
                END IF;

                IF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;

                b3 <= '1';

                b1 <= '0';

                b2 <= '1';

                b0 <= '1';
            WHEN ZE =>
                IF (NOT((x = '1'))) THEN
                    reg_fstate <= ZE;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= ZF;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= ZE;
                END IF;

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;

                b3 <= '1';

                b1 <= '1';

                b2 <= '1';

                b0 <= '0';
            WHEN ZF =>
                IF (NOT((x2 = '1'))) THEN
                    reg_fstate <= ZF;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= ZF;
                END IF;

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;

                b3 <= '1';

                b1 <= '1';

                b2 <= '1';

                b0 <= '1';
            WHEN vor =>
                IF ((x2 = '1')) THEN
                    reg_fstate <= vor2;
                ELSIF (NOT((x2 = '1'))) THEN
                    reg_fstate <= vor;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= vor;
                END IF;
            WHEN vor2 =>
                IF (NOT((x = '1'))) THEN
                    reg_fstate <= vor2;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= vor3;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= vor2;
                END IF;
            WHEN vor3 =>
                IF (NOT((x2 = '1'))) THEN
                    reg_fstate <= vor3;
                ELSIF ((x2 = '1')) THEN
                    reg_fstate <= Z0;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= vor3;
                END IF;
            WHEN OTHERS => 
                b3 <= 'X';
                b2 <= 'X';
                b1 <= 'X';
                b0 <= 'X';
                y <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
