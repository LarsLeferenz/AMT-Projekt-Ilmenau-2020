-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Wed Jun 24 18:37:12 2020

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY highacitve IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        x : IN STD_LOGIC := '0';
        y : OUT STD_LOGIC
    );
END highacitve;

ARCHITECTURE BEHAVIOR OF highacitve IS
    TYPE type_fstate IS (low,high,inactive);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= low;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,x)
    BEGIN
        y <= '0';
        CASE fstate IS
            WHEN low =>
                IF (NOT((x = '1'))) THEN
                    reg_fstate <= low;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= high;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= low;
                END IF;

                y <= '0';
            WHEN high =>
                IF ((x = '1')) THEN
                    reg_fstate <= inactive;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= high;
                END IF;

                y <= '1';
            WHEN inactive =>
                IF ((x = '1')) THEN
                    reg_fstate <= inactive;
                ELSIF (NOT((x = '1'))) THEN
                    reg_fstate <= low;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= inactive;
                END IF;

                y <= '0';
            WHEN OTHERS => 
                y <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
