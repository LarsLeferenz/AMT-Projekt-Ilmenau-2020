-- Copyright (C) 2019  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 19.1.0 Build 670 09/22/2019 SJ Lite Edition
-- Created on Mon Jul 27 11:55:43 2020

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY HEX_Counter IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        x : IN STD_LOGIC := '0';
        x2 : IN STD_LOGIC := '0';
        b3 : OUT STD_LOGIC;
        b2 : OUT STD_LOGIC;
        b1 : OUT STD_LOGIC;
        b0 : OUT STD_LOGIC;
        y : OUT STD_LOGIC
    );
END HEX_Counter;

ARCHITECTURE BEHAVIOR OF HEX_Counter IS
    TYPE type_fstate IS (Z0,Z1,Z2,Z3,Z4,Z5,Z6,Z7,Z8,Z9,ZA,ZB,ZC,ZD,ZE,ZF);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= Z0;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,x,x2)
    BEGIN
        b3 <= '0';
        b2 <= '0';
        b1 <= '0';
        b0 <= '0';
        y <= '0';
        CASE fstate IS
            WHEN Z0 =>
                IF (NOT((x = '1'))) THEN
                    reg_fstate <= Z0;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= Z1;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z0;
                END IF;

                b2 <= '0';

                b3 <= '0';

                b1 <= '0';

                b0 <= '0';

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;
                y <= '1';
            WHEN Z1 =>
                IF (NOT((x2 = '1'))) THEN
                    reg_fstate <= Z1;
                ELSIF ((x2 = '1')) THEN
                    reg_fstate <= Z2;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z1;
                END IF;

                b2 <= '0';

                b3 <= '0';

                b1 <= '0';

                b0 <= '1';

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;
            WHEN Z2 =>
                IF (NOT((x = '1'))) THEN
                    reg_fstate <= Z2;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= Z3;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z2;
                END IF;

                b2 <= '0';

                b3 <= '0';

                b1 <= '1';

                b0 <= '0';

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;
            WHEN Z3 =>
                IF (NOT((x2 = '1'))) THEN
                    reg_fstate <= Z3;
                ELSIF ((x2 = '1')) THEN
                    reg_fstate <= Z4;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z3;
                END IF;

                b2 <= '0';

                b3 <= '0';

                b1 <= '1';

                b0 <= '1';

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;
            WHEN Z4 =>
                IF (NOT((x = '1'))) THEN
                    reg_fstate <= Z4;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= Z5;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z4;
                END IF;

                b2 <= '1';

                b3 <= '0';

                b1 <= '0';

                b0 <= '0';

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;
            WHEN Z5 =>
                IF (NOT((x2 = '1'))) THEN
                    reg_fstate <= Z5;
                ELSIF ((x2 = '1')) THEN
                    reg_fstate <= Z6;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z5;
                END IF;

                b2 <= '1';

                b3 <= '0';

                b1 <= '0';

                b0 <= '1';

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;
            WHEN Z6 =>
                IF (NOT((x = '1'))) THEN
                    reg_fstate <= Z6;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= Z7;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z6;
                END IF;

                b2 <= '1';

                b3 <= '0';

                b1 <= '1';

                b0 <= '0';

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;
            WHEN Z7 =>
                IF (NOT((x2 = '1'))) THEN
                    reg_fstate <= Z7;
                ELSIF ((x2 = '1')) THEN
                    reg_fstate <= Z8;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z7;
                END IF;

                b2 <= '1';

                b3 <= '0';

                b1 <= '1';

                b0 <= '1';

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;
            WHEN Z8 =>
                IF (NOT((x = '1'))) THEN
                    reg_fstate <= Z8;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= Z9;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z8;
                END IF;

                b2 <= '0';

                b3 <= '1';

                b1 <= '0';

                b0 <= '0';

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;
            WHEN Z9 =>
                IF (NOT((x2 = '1'))) THEN
                    reg_fstate <= Z9;
                ELSIF ((x2 = '1')) THEN
                    reg_fstate <= ZA;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= Z9;
                END IF;

                b2 <= '0';

                b3 <= '1';

                b1 <= '0';

                b0 <= '1';

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;
            WHEN ZA =>
                IF (NOT((x = '1'))) THEN
                    reg_fstate <= ZA;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= ZB;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= ZA;
                END IF;

                b2 <= '0';

                b3 <= '1';

                b1 <= '1';

                b0 <= '0';

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;
            WHEN ZB =>
                IF (NOT((x2 = '1'))) THEN
                    reg_fstate <= ZB;
                ELSIF ((x2 = '1')) THEN
                    reg_fstate <= ZC;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= ZB;
                END IF;

                b2 <= '0';

                b3 <= '1';

                b1 <= '1';

                b0 <= '1';

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;
            WHEN ZC =>
                IF (NOT((x = '1'))) THEN
                    reg_fstate <= ZC;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= ZD;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= ZC;
                END IF;

                b2 <= '1';

                b3 <= '1';

                b1 <= '0';

                b0 <= '0';

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;
            WHEN ZD =>
                IF (NOT((x2 = '1'))) THEN
                    reg_fstate <= ZD;
                ELSIF ((x2 = '1')) THEN
                    reg_fstate <= ZE;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= ZD;
                END IF;

                b2 <= '1';

                b3 <= '1';

                b1 <= '0';

                b0 <= '1';

                IF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;
            WHEN ZE =>
                IF (NOT((x = '1'))) THEN
                    reg_fstate <= ZE;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= ZF;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= ZE;
                END IF;

                b2 <= '1';

                b3 <= '1';

                b1 <= '1';

                b0 <= '0';

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;
            WHEN ZF =>
                IF (NOT((x2 = '1'))) THEN
                    reg_fstate <= ZF;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= ZF;
                END IF;

                b2 <= '1';

                b3 <= '1';

                b1 <= '1';

                b0 <= '1';

                IF ((x = '1')) THEN
                    y <= '1';
                ELSIF (NOT((x = '1'))) THEN
                    y <= '0';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    y <= '0';
                END IF;
            WHEN OTHERS => 
                b3 <= 'X';
                b2 <= 'X';
                b1 <= 'X';
                b0 <= 'X';
                y <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
