// Copyright (C) 2019  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 19.1.0 Build 670 09/22/2019 SJ Lite Edition
// Created on Fri Aug 28 15:32:53 2020

// synthesis message_off 10175

`timescale 1ns/1ns

module pulsegenerator (
    clock,reset,x,
    y);

    input clock;
    input reset;
    input x;
    tri0 reset;
    tri0 x;
    output y;
    reg y;
    reg [2:0] fstate;
    reg [2:0] reg_fstate;
    parameter warten=0,set=1,warten2=2;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or x)
    begin
        if (reset) begin
            reg_fstate <= warten;
            y <= 1'b0;
        end
        else begin
            y <= 1'b0;
            case (fstate)
                warten: begin
                    if (x)
                        reg_fstate <= set;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= warten;

                    y <= 1'b0;
                end
                set: begin
                    reg_fstate <= warten2;

                    y <= 1'b1;
                end
                warten2: begin
                    if (~(x))
                        reg_fstate <= warten;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= warten2;

                    y <= 1'b0;
                end
                default: begin
                    y <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // pulsegenerator
