// Copyright (C) 2019  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 19.1.0 Build 670 09/22/2019 SJ Lite Edition
// Created on Mon Jul 20 16:37:07 2020

// synthesis message_off 10175

`timescale 1ns/1ns

module highacitve (
    clock,reset,x,
    y);

    input clock;
    input reset;
    input x;
    tri0 reset;
    tri0 x;
    output y;
    reg y;
    reg [2:0] fstate;
    reg [2:0] reg_fstate;
    parameter low=0,high=1,inactive=2;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or x)
    begin
        if (reset) begin
            reg_fstate <= low;
            y <= 1'b0;
        end
        else begin
            y <= 1'b0;
            case (fstate)
                low: begin
                    if (~(x))
                        reg_fstate <= low;
                    else if (x)
                        reg_fstate <= high;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= low;

                    y <= 1'b0;
                end
                high: begin
                    if (x)
                        reg_fstate <= inactive;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= high;

                    y <= 1'b1;
                end
                inactive: begin
                    if (x)
                        reg_fstate <= inactive;
                    else if (~(x))
                        reg_fstate <= low;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= inactive;

                    y <= 1'b0;
                end
                default: begin
                    y <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // highacitve
