-- Copyright (C) 2019  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 19.1.0 Build 670 09/22/2019 SJ Lite Edition
-- Created on Wed Jun 24 16:59:32 2020

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY takt_geber IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        SAL : IN STD_LOGIC := '0';
        stop : IN STD_LOGIC := '0';
        weiss : OUT STD_LOGIC;
        schwarz : OUT STD_LOGIC
    );
END takt_geber;

ARCHITECTURE BEHAVIOR OF takt_geber IS
    TYPE type_fstate IS (takt_wei�,takt_schwarz,halt);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= takt_wei�;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,SAL,stop)
    BEGIN
        weiss <= '0';
        schwarz <= '0';
        CASE fstate IS
            WHEN takt_wei� =>
                IF (((SAL = '1') AND NOT((stop = '1')))) THEN
                    reg_fstate <= takt_schwarz;
                ELSIF ((NOT((SAL = '1')) AND NOT((stop = '1')))) THEN
                    reg_fstate <= takt_wei�;
                ELSIF ((stop = '1')) THEN
                    reg_fstate <= halt;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= takt_wei�;
                END IF;

                weiss <= '1';

                schwarz <= '0';
            WHEN takt_schwarz =>
                IF ((NOT((SAL = '1')) AND NOT((stop = '1')))) THEN
                    reg_fstate <= takt_wei�;
                ELSIF (((SAL = '1') AND NOT((stop = '1')))) THEN
                    reg_fstate <= takt_schwarz;
                ELSIF ((stop = '1')) THEN
                    reg_fstate <= halt;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= takt_schwarz;
                END IF;

                weiss <= '0';

                schwarz <= '1';
            WHEN halt =>
                reg_fstate <= halt;
            WHEN OTHERS => 
                weiss <= 'X';
                schwarz <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
