-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Wed Jun 24 23:07:54 2020

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY d_flipflop IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        x : IN STD_LOGIC := '0';
        read : IN STD_LOGIC := '0';
        y : OUT STD_LOGIC
    );
END d_flipflop;

ARCHITECTURE BEHAVIOR OF d_flipflop IS
    TYPE type_fstate IS (one,zero);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x,read)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= zero;
            y <= '0';
        ELSE
            y <= '0';
            CASE fstate IS
                WHEN one =>
                    IF ((((x = '1') AND (read = '1')) OR NOT((read = '1')))) THEN
                        reg_fstate <= one;
                    ELSIF ((NOT((x = '1')) AND (read = '1'))) THEN
                        reg_fstate <= zero;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= one;
                    END IF;

                    y <= '1';
                WHEN zero =>
                    IF (((NOT((x = '1')) AND (read = '1')) OR NOT((read = '1')))) THEN
                        reg_fstate <= zero;
                    ELSIF (((x = '1') AND (read = '1'))) THEN
                        reg_fstate <= one;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= zero;
                    END IF;

                    y <= '0';
                WHEN OTHERS => 
                    y <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
