// Copyright (C) 2016  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Intel and sold by Intel or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// Generated by Quartus Prime Version 16.1.0 Build 196 10/24/2016 SJ Lite Edition
// Created on Mon Aug 14 15:11:45 2017

// synthesis message_off 10175

`timescale 1ns/1ns

module fahrstreckeVERILOG (reset,clock,fk,cl,cr,sl,sr,sk,dl,dr,ac,y3,y2,y1,y0);

    input reset;
    input clock;
    input fk;
	 input cl;
	 input cr;
	 
    tri0 reset;
    tri0 fk;
    tri0 cl;
    tri0 cr;
	 
    output sl;
    output sr;
    output sk;
    output dl;
    output dr;
	 output ac;
	 output y3;
    output y2;
    output y1;
    output y0;
    
    reg sl;
    reg sr;
    reg sk;
    reg dl;
    reg dr;
	 reg ac;
    reg y3;
    reg y2;
    reg y1;
    reg y0;
    
	 reg [4:0] fstate;
    reg [4:0] reg_fstate;
    parameter W1=0,W2=1,W3=2,W4=3,K1=4,K2=5,K3=6,Fertig=7;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or fk or cl or cr)
    begin
        if (~reset) begin
            reg_fstate <= W1;
            sl <= 1'b0;
            sr <= 1'b0;
            sk <= 1'b0;
            dl <= 1'b0;
            dr <= 1'b0;
				ac <= 1'b0;
        end
        else begin
            sl <= 1'b0;
            sr <= 1'b0;
            sk <= 1'b0;
            dl <= 1'b0;
            dr <= 1'b0;
            ac <= 1'b0;
				case (fstate)
					 W1: begin
                    if ((~(fk))&((~(cl))|(~(cr))))
                        reg_fstate <= W1;
                    else
                        reg_fstate <= K1;
                    // Inserting 'else' block to prevent latch inference

                    sk <= 1'b0;

                    sr <= 1'b0;

                    sl <= 1'b0;

                    dr <= 1'b0;

                    dl <= 1'b0;
						  
						  ac <= 1'b0;
						  
						  y3 <= 0;
						  y2 <= 0;
						  y1 <= 0;
						  y0 <= 0; 
                end
                K1: begin
                    if ((~(fk))&((~(cl))|(~(cr))))
                        reg_fstate <= W2;
                    else
								reg_fstate <= K1;
                    // Inserting 'else' block to prevent latch inference


                    sk <= 1'b0;

                    sr <= 1'b1;

                    sl <= 1'b0;

                    dr <= 1'b0;

                    dl <= 1'b0;
						  
						  ac <= 1'b1;
						  
						  y3 <= 0;
						  y2 <= 0;
						  y1 <= 0;
						  y0 <= 1; 
                end
                
					 W2: begin
                    if ((~(fk))&((~(cl))|(~(cr))))
                        reg_fstate <= W2;
                    else
                        reg_fstate <= K2;
                    // Inserting 'else' block to prevent latch inference

                    sk <= 1'b0;

                    sr <= 1'b0;

                    sl <= 1'b0;

                    dr <= 1'b0;

                    dl <= 1'b0;
						  
						  ac <= 1'b0;
						  
						  y3 <= 0;
						  y2 <= 0;
						  y1 <= 1;
						  y0 <= 0; 
                end
                K2: begin
                    if ((~(fk))&((~(cl))|(~(cr))))
                        reg_fstate <= W3;
                    else
								reg_fstate <= K2;
                    // Inserting 'else' block to prevent latch inference


                    sk <= 1'b1;

                    sr <= 1'b0;

                    sl <= 1'b0;

                    dr <= 1'b0;

                    dl <= 1'b0;
						  
						  ac <= 1'b1;
						  
						  y3 <= 0;
						  y2 <= 0;
						  y1 <= 1;
						  y0 <= 1; 
                end
					 
					 W3: begin
                    if ((~(fk))&((~(cl))|(~(cr))))
                        reg_fstate <= W3;
                    else
                        reg_fstate <= K3;
                    // Inserting 'else' block to prevent latch inference

                    sk <= 1'b0;

                    sr <= 1'b0;

                    sl <= 1'b0;

                    dr <= 1'b0;

                    dl <= 1'b0;
						  
						  ac <= 1'b1;
						  
						  y3 <= 0;
						  y2 <= 1;
						  y1 <= 0;
						  y0 <= 0; 
                end
                K3: begin
                    if ((~(fk))&((~(cl))|(~(cr))))
                        reg_fstate <= W4;
                    else
								reg_fstate <= K3;
                    // Inserting 'else' block to prevent latch inference


                    sk <= 1'b0;

                    sr <= 1'b1;

                    sl <= 1'b0;

                    dr <= 1'b0;

                    dl <= 1'b0;
						  
						  ac <= 1'b0;
						  
						  y3 <= 0;
						  y2 <= 1;
						  y1 <= 0;
						  y0 <= 1; 
                end
					 
					 W4: begin
                    if ((~(fk))&((~(cl))|(~(cr))))
                        reg_fstate <= W4;
                    else
                        reg_fstate <= Fertig;
                    // Inserting 'else' block to prevent latch inference

                    sk <= 1'b0;

                    sr <= 1'b0;

                    sl <= 1'b0;

                    dr <= 1'b0;

                    dl <= 1'b0;
						  
						  ac <= 1'b1;
						  
						  y3 <= 0;
						  y2 <= 1;
						  y1 <= 1;
						  y0 <= 0; 
                end
                
                Fertig: begin
                    reg_fstate <= Fertig;

                    sk <= 1'b0;

                    sr <= 1'b0;

                    sl <= 1'b0;

                    dr <= 1'b0;

                    dl <= 1'b1;
						  
						  ac <= 1'b1;
						  
						  y3 <= 0;
						  y2 <= 1;
						  y1 <= 1;
						  y0 <= 1; 
                end
                default: begin
                    sl <= 1'bx;
                    sr <= 1'bx;
                    sk <= 1'bx;
                    dl <= 1'bx;
                    dr <= 1'bx;
						  ac <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // fahrstrecke
