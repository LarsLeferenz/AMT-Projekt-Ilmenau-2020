-- Copyright (C) 2016  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Intel and sold by Intel or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- Generated by Quartus Prime Version 16.1.0 Build 196 10/24/2016 SJ Lite Edition
-- Created on Tue Sep 05 13:39:41 2017

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY fahrsteuerung IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        xkl : IN STD_LOGIC := '0';
        xkr : IN STD_LOGIC := '0';
        xll : IN STD_LOGIC := '0';
        xlr : IN STD_LOGIC := '0';
        sl : IN STD_LOGIC := '0';
        sr : IN STD_LOGIC := '0';
        dl : IN STD_LOGIC := '0';
        dr : IN STD_LOGIC := '0';
        ac : IN STD_LOGIC := '0';
        delayReady : IN STD_LOGIC := '0';
        ready : IN STD_LOGIC := '0';
        stop : IN STD_LOGIC := '0';
        yml : OUT STD_LOGIC;
        ymr : OUT STD_LOGIC;
        ymlr : OUT STD_LOGIC;
        ymrr : OUT STD_LOGIC;
        cl : OUT STD_LOGIC;
        cr : OUT STD_LOGIC;
        fk : OUT STD_LOGIC;
        z0 : OUT STD_LOGIC;
        z1 : OUT STD_LOGIC;
        z2 : OUT STD_LOGIC;
        delayStart : OUT STD_LOGIC;
        z3 : OUT STD_LOGIC
    );
END fahrsteuerung;

ARCHITECTURE BEHAVIOR OF fahrsteuerung IS
    TYPE type_fstate IS (IdleFahren,Abzweig,LinieRechts,KurveRechts,LinieLinks,KurveLinks,KreiselnRechts,KreiselnLinks,WarteLinks,DreheLinks,WarteRechts,DreheRechts,WarteAufLinieLinks,WarteAufLinieRechts);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,xkl,xkr,xll,xlr,sl,sr,dl,dr,ac,delayReady,ready,stop)
    BEGIN
        IF (reset='0') THEN
            reg_fstate <= IdleFahren;
            yml <= '0';
            ymr <= '0';
            ymlr <= '0';
            ymrr <= '0';
            cl <= '0';
            cr <= '0';
            fk <= '0';
            z0 <= '0';
            z1 <= '0';
            z2 <= '0';
            delayStart <= '0';
            z3 <= '0';
        ELSE
            yml <= '0';
            ymr <= '0';
            ymlr <= '0';
            ymrr <= '0';
            cl <= '0';
            cr <= '0';
            fk <= '0';
            z0 <= '0';
            z1 <= '0';
            z2 <= '0';
            delayStart <= '0';
            z3 <= '0';
            CASE fstate IS
                WHEN IdleFahren =>
                    IF (((ready = '1') AND ((((xkr = '1') AND NOT((dr = '1'))) AND NOT((dl = '1'))) OR (((xkl = '1') AND NOT((dr = '1'))) AND NOT((dl = '1')))))) THEN
                        reg_fstate <= Abzweig;
                    ELSIF ((((dr = '1') AND NOT((dl = '1'))) AND (ready = '1'))) THEN
                        reg_fstate <= KreiselnRechts;
                    ELSIF (((NOT((dr = '1')) AND (dl = '1')) AND (ready = '1'))) THEN
                        reg_fstate <= KreiselnLinks;
                    ELSIF ((((((NOT((xkr = '1')) AND NOT((xkl = '1'))) AND NOT((dr = '1'))) AND NOT((dl = '1'))) OR ((dl = '1') AND (dr = '1'))) OR NOT((ready = '1')))) THEN
                        reg_fstate <= IdleFahren;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= IdleFahren;
                    END IF;

                    z3 <= '0';

                    z2 <= '0';

                    z1 <= '0';

                    z0 <= '0';

                    fk <= '0';

                    cr <= '0';

                    cl <= '0';

                    ymrr <= '0';

                    ymlr <= '0';

                    ymr <= (xll AND NOT(stop));

                    yml <= (xlr AND NOT(stop));

                    delayStart <= '0';
                WHEN Abzweig =>
                    IF ((NOT((xkr = '1')) AND NOT((xkl = '1')))) THEN
                        reg_fstate <= IdleFahren;
                    ELSIF (((((xkr = '1') AND (sr = '1')) AND NOT((sl = '1'))) AND NOT((ac = '1')))) THEN
                        reg_fstate <= KurveRechts;
                    ELSIF (((((xkl = '1') AND NOT((sr = '1'))) AND (sl = '1')) AND NOT((ac = '1')))) THEN
                        reg_fstate <= KurveLinks;
                    ELSIF (((((xkl = '1') AND NOT((sr = '1'))) AND (sl = '1')) AND (ac = '1'))) THEN
                        reg_fstate <= WarteLinks;
                    ELSIF (((((xkr = '1') AND (sr = '1')) AND NOT((sl = '1'))) AND (ac = '1'))) THEN
                        reg_fstate <= WarteRechts;
                    ELSIF (((((((xkl = '1') AND NOT((sl = '1'))) AND NOT((sr = '1'))) OR (((xkr = '1') AND NOT((xkl = '1'))) AND NOT((sr = '1')))) OR (((xkr = '1') AND (sr = '1')) AND (sl = '1'))) OR ((NOT((xkr = '1')) AND (xkl = '1')) AND (sr = '1')))) THEN
                        reg_fstate <= Abzweig;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Abzweig;
                    END IF;

                    z3 <= '0';

                    z2 <= '0';

                    z1 <= '0';

                    z0 <= '1';

                    fk <= '0';

                    cr <= xkr;

                    cl <= xkl;

                    ymrr <= '0';

                    ymlr <= '0';

                    ymr <= ((((xkl AND NOT((sr AND sl))) OR (xkl AND sl)) OR (NOT(xlr) AND xkr)) AND NOT(stop));

                    yml <= ((((xkr AND NOT((sr AND sl))) OR (xkr AND sr)) OR (NOT(xll) AND xkl)) AND NOT(stop));

                    delayStart <= '0';
                WHEN LinieRechts =>
                    IF ((xll = '1')) THEN
                        reg_fstate <= IdleFahren;
                    ELSIF (NOT((xll = '1'))) THEN
                        reg_fstate <= LinieRechts;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= LinieRechts;
                    END IF;

                    z3 <= '0';

                    z2 <= '0';

                    z1 <= '1';

                    z0 <= '0';

                    fk <= '1';

                    cr <= '0';

                    cl <= '0';

                    ymrr <= '0';

                    ymlr <= '0';

                    ymr <= '0';

                    yml <= NOT(stop);

                    delayStart <= '0';
                WHEN KurveRechts =>
                    IF (NOT((xll = '1'))) THEN
                        reg_fstate <= LinieRechts;
                    ELSIF ((xll = '1')) THEN
                        reg_fstate <= KurveRechts;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= KurveRechts;
                    END IF;

                    z3 <= '0';

                    z2 <= '0';

                    z1 <= '1';

                    z0 <= '1';

                    fk <= '1';

                    cr <= '0';

                    cl <= '0';

                    ymrr <= '0';

                    ymlr <= '0';

                    ymr <= '0';

                    yml <= NOT(stop);

                    delayStart <= '0';
                WHEN LinieLinks =>
                    IF ((xlr = '1')) THEN
                        reg_fstate <= IdleFahren;
                    ELSIF (NOT((xlr = '1'))) THEN
                        reg_fstate <= LinieLinks;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= LinieLinks;
                    END IF;

                    z3 <= '0';

                    z2 <= '1';

                    z1 <= '0';

                    z0 <= '0';

                    fk <= '1';

                    cr <= '0';

                    cl <= '0';

                    ymrr <= '0';

                    ymlr <= '0';

                    ymr <= NOT(stop);

                    yml <= '0';

                    delayStart <= '0';
                WHEN KurveLinks =>
                    IF (NOT((xlr = '1'))) THEN
                        reg_fstate <= LinieLinks;
                    ELSIF ((xlr = '1')) THEN
                        reg_fstate <= KurveLinks;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= KurveLinks;
                    END IF;

                    z3 <= '0';

                    z2 <= '1';

                    z1 <= '0';

                    z0 <= '1';

                    fk <= '1';

                    cr <= '0';

                    cl <= '0';

                    ymrr <= '0';

                    ymlr <= '0';

                    ymr <= NOT(stop);

                    yml <= '0';

                    delayStart <= '0';
                WHEN KreiselnRechts =>
                    reg_fstate <= KreiselnRechts;

                    z3 <= '1';

                    z2 <= '1';

                    z1 <= '0';

                    z0 <= '0';

                    fk <= '0';

                    cr <= '0';

                    cl <= '0';

                    ymrr <= '1';

                    ymlr <= '0';

                    ymr <= '0';

                    yml <= '1';

                    delayStart <= '0';
                WHEN KreiselnLinks =>
                    reg_fstate <= KreiselnLinks;

                    z3 <= '1';

                    z2 <= '1';

                    z1 <= '0';

                    z0 <= '1';

                    fk <= '0';

                    cr <= '0';

                    cl <= '0';

                    ymrr <= '0';

                    ymlr <= NOT(stop);

                    ymr <= '1';

                    yml <= '0';

                    delayStart <= '0';
                WHEN WarteLinks =>
                    IF ((delayReady = '1')) THEN
                        reg_fstate <= DreheLinks;
                    ELSIF (NOT((delayReady = '1'))) THEN
                        reg_fstate <= WarteLinks;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= WarteLinks;
                    END IF;

                    z3 <= '1';

                    z2 <= '0';

                    z1 <= '0';

                    z0 <= '0';

                    fk <= '1';

                    cr <= '0';

                    cl <= '0';

                    ymrr <= '0';

                    ymlr <= '0';

                    ymr <= NOT(stop);

                    yml <= NOT(stop);

                    delayStart <= '1';
                WHEN DreheLinks =>
                    IF ((NOT((xlr = '1')) AND NOT((xll = '1')))) THEN
                        reg_fstate <= WarteAufLinieLinks;
                    ELSIF (((xlr = '1') OR (xll = '1'))) THEN
                        reg_fstate <= DreheLinks;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= DreheLinks;
                    END IF;

                    z3 <= '1';

                    z2 <= '0';

                    z1 <= '0';

                    z0 <= '1';

                    fk <= '1';

                    cr <= '0';

                    cl <= '0';

                    ymrr <= '0';

                    ymlr <= NOT(stop);

                    ymr <= NOT(stop);

                    yml <= '0';

                    delayStart <= '0';
                WHEN WarteRechts =>
                    IF ((delayReady = '1')) THEN
                        reg_fstate <= DreheRechts;
                    ELSIF (NOT((delayReady = '1'))) THEN
                        reg_fstate <= WarteRechts;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= WarteRechts;
                    END IF;

                    z3 <= '0';

                    z2 <= '1';

                    z1 <= '1';

                    z0 <= '0';

                    fk <= '1';

                    cr <= '0';

                    cl <= '0';

                    ymrr <= '0';

                    ymlr <= '0';

                    ymr <= NOT(stop);

                    yml <= NOT(stop);

                    delayStart <= '1';
                WHEN DreheRechts =>
                    IF ((NOT((xll = '1')) AND NOT((xlr = '1')))) THEN
                        reg_fstate <= WarteAufLinieRechts;
                    ELSIF (((xll = '1') OR (xlr = '1'))) THEN
                        reg_fstate <= DreheRechts;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= DreheRechts;
                    END IF;

                    z3 <= '0';

                    z2 <= '1';

                    z1 <= '1';

                    z0 <= '1';

                    fk <= '1';

                    cr <= '0';

                    cl <= '0';

                    ymrr <= NOT(stop);

                    ymlr <= '0';

                    ymr <= '0';

                    yml <= NOT(stop);

                    delayStart <= '0';
                WHEN WarteAufLinieLinks =>
                    IF ((xlr = '1')) THEN
                        reg_fstate <= IdleFahren;
                    ELSIF (NOT((xlr = '1'))) THEN
                        reg_fstate <= WarteAufLinieLinks;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= WarteAufLinieLinks;
                    END IF;

                    z3 <= '1';

                    z2 <= '0';

                    z1 <= '1';

                    z0 <= '1';

                    fk <= '1';

                    cr <= '0';

                    cl <= '0';

                    ymrr <= '0';

                    ymlr <= NOT(stop);

                    ymr <= NOT(stop);

                    yml <= '0';

                    delayStart <= '0';
                WHEN WarteAufLinieRechts =>
                    IF ((xll = '1')) THEN
                        reg_fstate <= IdleFahren;
                    ELSIF (NOT((xll = '1'))) THEN
                        reg_fstate <= WarteAufLinieRechts;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= WarteAufLinieRechts;
                    END IF;

                    z3 <= '1';

                    z2 <= '0';

                    z1 <= '1';

                    z0 <= '0';

                    fk <= '1';

                    cr <= '0';

                    cl <= '0';

                    ymrr <= NOT(stop);

                    ymlr <= '0';

                    ymr <= '0';

                    yml <= NOT(stop);

                    delayStart <= '0';
                WHEN OTHERS => 
                    yml <= 'X';
                    ymr <= 'X';
                    ymlr <= 'X';
                    ymrr <= 'X';
                    cl <= 'X';
                    cr <= 'X';
                    fk <= 'X';
                    z0 <= 'X';
                    z1 <= 'X';
                    z2 <= 'X';
                    delayStart <= 'X';
                    z3 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
