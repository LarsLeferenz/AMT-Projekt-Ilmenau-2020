-- Copyright (C) 2019  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 19.1.0 Build 670 09/22/2019 SJ Lite Edition
-- Created on Fri Aug 28 18:07:18 2020

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY NFolge IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        sli : IN STD_LOGIC := '0';
        sri : IN STD_LOGIC := '0';
        sar : IN STD_LOGIC := '0';
        sal : IN STD_LOGIC := '0';
        y0 : IN STD_LOGIC := '0';
        y1 : IN STD_LOGIC := '0';
        mlv : OUT STD_LOGIC;
        mrv : OUT STD_LOGIC;
        mlr : OUT STD_LOGIC;
        mrr : OUT STD_LOGIC;
        Kreuzung : OUT STD_LOGIC
    );
END NFolge;

ARCHITECTURE BEHAVIOR OF NFolge IS
    TYPE type_fstate IS (gerade,links,rechts,kreuz,kreuzab,schlinks,schrechts,kreuzauf,kreuzlink,kreuzrech,KreuzLeer);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,sli,sri,sar,sal,y0,y1)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= gerade;
            mlv <= '0';
            mrv <= '0';
            mlr <= '0';
            mrr <= '0';
            Kreuzung <= '0';
        ELSE
            mlv <= '0';
            mrv <= '0';
            mlr <= '0';
            mrr <= '0';
            Kreuzung <= '0';
            CASE fstate IS
                WHEN gerade =>
                    IF (((((sli = '1') AND (sri = '1')) AND NOT((sal = '1'))) AND NOT((sar = '1')))) THEN
                        reg_fstate <= gerade;
                    ELSIF (((((sli = '1') AND NOT((sri = '1'))) AND NOT((sal = '1'))) AND NOT((sar = '1')))) THEN
                        reg_fstate <= links;
                    ELSIF ((((NOT((sli = '1')) AND (sri = '1')) AND NOT((sal = '1'))) AND NOT((sar = '1')))) THEN
                        reg_fstate <= rechts;
                    ELSIF ((((sli = '1') OR (sri = '1')) AND ((sal = '1') OR (sar = '1')))) THEN
                        reg_fstate <= kreuzauf;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= gerade;
                    END IF;

                    mlr <= '0';

                    mrr <= '0';

                    mlv <= '1';

                    mrv <= '1';

                    Kreuzung <= '0';
                WHEN links =>
                    IF (((sli = '1') AND NOT((sri = '1')))) THEN
                        reg_fstate <= links;
                    ELSIF ((sri = '1')) THEN
                        reg_fstate <= gerade;
                    ELSIF ((NOT((sli = '1')) AND NOT((sri = '1')))) THEN
                        reg_fstate <= schlinks;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= links;
                    END IF;

                    mlr <= '0';

                    mrr <= '0';

                    mlv <= '0';

                    mrv <= '1';

                    Kreuzung <= '0';
                WHEN rechts =>
                    IF ((NOT((sli = '1')) AND (sri = '1'))) THEN
                        reg_fstate <= rechts;
                    ELSIF ((sli = '1')) THEN
                        reg_fstate <= gerade;
                    ELSIF ((NOT((sli = '1')) AND NOT((sri = '1')))) THEN
                        reg_fstate <= schrechts;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= rechts;
                    END IF;

                    mlr <= '0';

                    mrr <= '0';

                    mlv <= '1';

                    mrv <= '0';

                    Kreuzung <= '0';
                WHEN kreuz =>
                    IF ((NOT((sal = '1')) AND NOT((sar = '1')))) THEN
                        reg_fstate <= kreuzab;
                    ELSIF (((sal = '1') OR (sar = '1'))) THEN
                        reg_fstate <= kreuz;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= kreuz;
                    END IF;

                    mlr <= '0';

                    mrr <= '0';

                    mlv <= '1';

                    mrv <= '1';

                    Kreuzung <= '0';
                WHEN kreuzab =>
                    reg_fstate <= gerade;

                    mlr <= '0';

                    mrr <= '0';

                    mlv <= '0';

                    mrv <= '0';

                    Kreuzung <= '1';
                WHEN schlinks =>
                    IF (NOT((sli = '1'))) THEN
                        reg_fstate <= schlinks;
                    ELSIF ((sli = '1')) THEN
                        reg_fstate <= links;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= schlinks;
                    END IF;

                    mlr <= '1';

                    mrr <= '0';

                    mlv <= '0';

                    mrv <= '1';

                    Kreuzung <= '0';
                WHEN schrechts =>
                    IF (NOT((sri = '1'))) THEN
                        reg_fstate <= schrechts;
                    ELSIF ((sri = '1')) THEN
                        reg_fstate <= rechts;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= schrechts;
                    END IF;

                    mlr <= '0';

                    mrr <= '1';

                    mlv <= '1';

                    mrv <= '0';

                    Kreuzung <= '0';
                WHEN kreuzauf =>
                    IF ((NOT((y0 = '1')) AND (y1 = '1'))) THEN
                        reg_fstate <= kreuzlink;
                    ELSIF (((y0 = '1') AND (y1 = '1'))) THEN
                        reg_fstate <= kreuz;
                    ELSIF (((y0 = '1') AND NOT((y1 = '1')))) THEN
                        reg_fstate <= kreuzrech;
                    ELSIF ((NOT((y0 = '1')) AND NOT((y1 = '1')))) THEN
                        reg_fstate <= KreuzLeer;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= kreuzauf;
                    END IF;

                    mlr <= '0';

                    mrr <= '0';

                    mlv <= '1';

                    mrv <= '1';

                    Kreuzung <= '0';
                WHEN kreuzlink =>
                    IF ((sri = '1')) THEN
                        reg_fstate <= kreuzlink;
                    ELSIF (NOT((sri = '1'))) THEN
                        reg_fstate <= links;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= kreuzlink;
                    END IF;

                    mlr <= '0';

                    mrr <= '0';

                    mlv <= '0';

                    mrv <= '1';

                    Kreuzung <= '1';
                WHEN kreuzrech =>
                    IF ((sli = '1')) THEN
                        reg_fstate <= kreuzrech;
                    ELSIF (NOT((sli = '1'))) THEN
                        reg_fstate <= rechts;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= kreuzrech;
                    END IF;

                    mlr <= '0';

                    mrr <= '0';

                    mlv <= '1';

                    mrv <= '0';

                    Kreuzung <= '1';
                WHEN KreuzLeer =>
                    reg_fstate <= kreuz;
                WHEN OTHERS => 
                    mlv <= 'X';
                    mrv <= 'X';
                    mlr <= 'X';
                    mrr <= 'X';
                    Kreuzung <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
