-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Fri Aug 28 15:37:39 2020

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY flipflop IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        x : IN STD_LOGIC := '0';
        y1 : OUT STD_LOGIC;
        y2 : OUT STD_LOGIC
    );
END flipflop;

ARCHITECTURE BEHAVIOR OF flipflop IS
    TYPE type_fstate IS (wait1,active1,wait2,active2);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= wait1;
            y1 <= '0';
            y2 <= '0';
        ELSE
            y1 <= '0';
            y2 <= '0';
            CASE fstate IS
                WHEN wait1 =>
                    IF (NOT((x = '1'))) THEN
                        reg_fstate <= wait1;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= active1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= wait1;
                    END IF;

                    y2 <= '1';

                    y1 <= '0';
                WHEN active1 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= active1;
                    ELSIF (NOT((x = '1'))) THEN
                        reg_fstate <= wait2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= active1;
                    END IF;

                    y2 <= '0';

                    y1 <= '1';
                WHEN wait2 =>
                    IF (NOT((x = '1'))) THEN
                        reg_fstate <= wait2;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= active2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= wait2;
                    END IF;

                    y2 <= '0';

                    y1 <= '1';
                WHEN active2 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= active2;
                    ELSIF (NOT((x = '1'))) THEN
                        reg_fstate <= wait1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= active2;
                    END IF;

                    y2 <= '1';

                    y1 <= '0';
                WHEN OTHERS => 
                    y1 <= 'X';
                    y2 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
