-- Copyright (C) 2019  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 19.1.0 Build 670 09/22/2019 SJ Lite Edition
-- Created on Wed Jun 24 16:46:00 2020

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY einlese_automat IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        schwarz : IN STD_LOGIC := '0';
        weiss : IN STD_LOGIC := '0';
        SAR : IN STD_LOGIC := '0';
        s0 : OUT STD_LOGIC;
        s1 : OUT STD_LOGIC;
        lesen : OUT STD_LOGIC
    );
END einlese_automat;

ARCHITECTURE BEHAVIOR OF einlese_automat IS
    TYPE type_fstate IS (start,erstes_schwarz,erstes_wei�,zweites_schwarz,zweites_wei�,erstes_schwarz_warten,erstes_wei�_warten);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= start;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,schwarz,weiss,SAR)
    BEGIN
        s0 <= '0';
        s1 <= '0';
        lesen <= '0';
        CASE fstate IS
            WHEN start =>
                IF (((SAR = '1') AND (weiss = '1'))) THEN
                    reg_fstate <= erstes_schwarz;
                ELSIF ((NOT((SAR = '1')) AND (weiss = '1'))) THEN
                    reg_fstate <= erstes_wei�;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= start;
                END IF;

                lesen <= '0';

                s1 <= '0';

                s0 <= '0';
            WHEN erstes_schwarz =>
                IF ((schwarz = '1')) THEN
                    reg_fstate <= erstes_schwarz_warten;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= erstes_schwarz;
                END IF;

                s0 <= '1';
            WHEN erstes_wei� =>
                IF ((schwarz = '1')) THEN
                    reg_fstate <= erstes_wei�_warten;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= erstes_wei�;
                END IF;
            WHEN zweites_schwarz =>
                IF ((schwarz = '1')) THEN
                    reg_fstate <= start;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= zweites_schwarz;
                END IF;

                lesen <= '1';

                s1 <= '1';
            WHEN zweites_wei� =>
                IF ((schwarz = '1')) THEN
                    reg_fstate <= start;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= zweites_wei�;
                END IF;

                lesen <= '1';
            WHEN erstes_schwarz_warten =>
                IF (((SAR = '1') AND (weiss = '1'))) THEN
                    reg_fstate <= zweites_schwarz;
                ELSIF ((NOT((SAR = '1')) AND (weiss = '1'))) THEN
                    reg_fstate <= zweites_wei�;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= erstes_schwarz_warten;
                END IF;
            WHEN erstes_wei�_warten =>
                IF (((SAR = '1') AND (weiss = '1'))) THEN
                    reg_fstate <= zweites_schwarz;
                ELSIF ((NOT((SAR = '1')) AND (weiss = '1'))) THEN
                    reg_fstate <= zweites_wei�;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= erstes_wei�_warten;
                END IF;
            WHEN OTHERS => 
                s0 <= 'X';
                s1 <= 'X';
                lesen <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
